/*
 * Copyright (c) 2025 Bennett Miller
 * SPDX-License-Identifier: Apache-2.0
 */

module tt_um_big_ben_fr_implies_gate (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // first four bits -> A, next four bits -> B

  wire [3:0] A = ui_in[3:0];
  wire [3:0] B = ui_in[7:4];

  assign uo_out[3:0] = ~(A) | B;

  assign uo_out[7:4] = 0; 
  assign uio_out = 0;
  assign uio_oe  = 0;

  wire _unused = &{ena, clk, rst_n, 1'b0};

endmodule